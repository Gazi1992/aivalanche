
.subckt dut p n

******* Junction DC parameters
+ IS=1e-14 JSW=1e-15 N=1 RS=0 BV=1e10 IBV=1e-3 NBV=1 IKF=0 IKR=0
+ JTUN=0 JTUNSW=0 NTUN=30 XTITUN=3 KEG=1 ISR=1e-14 NR=1

******* Junction capacitance parameters
+ CJO=0 CJP=0 FC=0.5 FCS=0.5 M=0.5 MJSW=0.33 VJ=1 PHP=1 TT=0

******* Metal and Polysilicon Overlap Capacitances (level=3)
+ LM=0 LP=0 WM=0 WP=0 XOM=1e-6 XOI=1e-6 XM=0 XP=0

******* Temperature effects
+ EG=1.11 TNOM=27 TRS1=0 TRS2=0 TM1=0 TM2=0 TTT1=0 TTT2=0 XTI=3
+ TLEV=0 TLEVC=0 CTA=0 CTP=0 TCV=0

******* Noise modeling
+ KF=0 AF=1


.model diode D

******* Junction DC parameters
+ IS=IS JSW=JSW N=N RS=RS BV=BV IBV=IBV NBV=NBV IKF=IKF IKR=IKR
+ JTUN=JTUN JTUNSW=JTUNSW NTUN=NTUN XTITUN=XTITUN KEG=KEG ISR=ISR NR=NR

******* Junction capacitance parameters
+ CJO=CJO CJP=CJP FC=FC FCS=FCS M=M MJSW=MJSW VJ=VJ PHP=PHP TT=TT

******* Metal and Polysilicon Overlap Capacitances (level=3)
+ LM=LM LP=LP WM=WM WP=WP XOM=XOM XOI=XOI XM=XM XP=XP

******* Temperature effects
+ EG=EG TNOM=TNOM TRS1=TRS1 TRS2=TRS2 TM1=TM1 TM2=TM2 TTT1=TTT1 TTT2=TTT2 XTI=XTI
+ TLEV=TLEV TLEVC=TLEVC CTA=CTA CTP=CTP TCV=TCV

******* Noise modeling
+ KF=KF AF=AF


d1 p n diode

.ends
