
.include dut1.cir

******************************* dut testbench 1 *******************************
vgs_1_ac g_1 g_1_ac DC 0 AC 1
egs_1 g_1_ac 0 v_sweep 0 1
vds_1 d_1 0 0
vs_1 s_1 0 0
vbs_1 b_1 0 0
x_1 d_1 g_1 s_1 b_1 dut l=5e-6 w=10e-1
*******************************************************************************

v_sweep v_sweep 0 DC 0

******************************* save data to file *****************************
.control

echo "v(g_1),cgd,cgs,cgb,cgg" > cgg_characteristic_results.csv

** Start the simulation loop.
*set values_list = ( 0.0 0.2 0.3 0.4 0.5 0.6 0.7 0.8 0.9 1.0 1.1 1.2 1.3 1.4 1.5 1.6 )
compose values_list start=-0.5 stop=3.5 step=0.05
print values_list
let kot = unitvec(length(values_list))
let i = 0

foreach val $&values_list

alter v_sweep $val
ac lin 3 1k 10k

let temp_cgg = (abs(imag(i(vds_1))) + abs(imag(i(vbs_1))) + abs(imag(i(vs_1))))/2*pi*10000
let temp_cgd = abs(imag(i(vds_1)))/2*pi*10000
let temp_cgs = abs(imag(i(vs_1)))/2*pi*10000
let temp_cgb = abs(imag(i(vbs_1)))/2*pi*10000

meas AC cgg FIND temp_cgg AT=10k
meas AC cgd FIND temp_cgd AT=10k
meas AC cgs FIND temp_cgs AT=10k
meas AC cgb FIND temp_cgb AT=10k

echo "$val,$&cgd,$&cgs,$&cgb,$&cgg" >> cgg_characteristic_results.csv

let i = i + 1
let kot[i] = cgg
end

.endc
*******************************************************************************

.end