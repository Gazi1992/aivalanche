** Single NMOS Transistor .measure (Id-Vd) **
* Altering device width leads to select new model due to binning limits.
* New model has artificially thick gate oxide (changed from default 3n to 4n)
* to demonstrate the effect.

* model binning
* uses default parameters, except toxe
* level 54 specifies the BSIM4 model
.model nch nmos level=54

m1 d g s b nch L=5e-6 W=10e-6  

vgs g 0 3.5
vds d 0 3.5
vs s 0 dc 0
vb b 0 dc 0

.control
dc vds 0 3.5 0.05 vgs 3.5 0.5 -0.5
set wr_vecnames
set wr_singlescale
wrdata Result.txt i(vs) v(d) v(g)
.endc

.end