
.include dut1.cir

******************************* dut testbench 1 *******************************
vgs_ac_1 g_1 g_1_ac DC 0 AC 1
egs_1 g_1_ac 0 v_sweep 0 1
vds_1 d_1 0 0
vs_1 s_1 0 0
vbs_1 b_1 0 0
x_1 d_1 g_1 s_1 b_1 dut l=5e-6 w=10e-1
*******************************************************************************

v_sweep v_sweep 0 DC 0

******************************* save data to file *****************************
.control

echo "v(g_1),cgd,cgs,cgb,cgg" > cgg_characteristic_results.csv

** Start the simulation loop.
compose values_list start=-0.5 stop=3.5 step=0.05
foreach val $&values_list
    alter v_sweep $val
    ac lin 1 10k 10k
    
    let cgd = abs(imag(i(vds_1)))/2*pi*10000
    let cgs = abs(imag(i(vs_1)))/2*pi*10000
    let cgb = abs(imag(i(vbs_1)))/2*pi*10000
    let cgg = (abs(imag(i(vds_1))) + abs(imag(i(vbs_1))) + abs(imag(i(vs_1))))/2*pi*10000
 
    echo "$val,$&cgd,$&cgs,$&cgb,$&cgg" >> cgg_characteristic_results.csv
end

.endc
*******************************************************************************

.end