
.subckt dut d g s b
* instance parameters
+ l = 10e-6
+ w = 10e-6
* model parameters
+ vth0 = 0.5
+ TNOM = 27


.model nch nmos version=4.8 level=54
* instance parameters
+ l = l
+ w = w
* model parameters
+ vth0 = vth0
+ TNOM = TNOM


m1 d g s b nch

.ends
