********** BSIM4 NMOS TEMPLATE **********

.subckt dut d g s b
********** instance parameters **********
+ l = 10e-6
+ w = 10e-6
+ nf = 1
+ m = 1
+ sa = 0
+ sb = 0
+ sc = 0
+ sca = 1
+ scb = 1
+ scc = 1
+ ad = 1e-12
+ pd = 1e-6
+ as = 1e-12
+ ps = 1e-6
+ nrs = 1
+ nrd = 1
********** model parameters **********
+ binunit = 1
+ paramchk = 0
+ mobmod = 0
+ capmod = 2
+ rdsmod = 0
+ igcmod = 0
+ igbmod = 0
+ rbodymod = 0
+ trnqsmod = 0
+ acnqsmod = 0
+ fnoimod = 1
+ tnoimod = 0
+ diomod = 1
+ tempmod = 2
+ permod = 1
+ geomod = 0
+ rgeomod = 0
+ rgatemod = 0
+ wpemod = 0
+ lmax = 1E-4
+ wmax = 1
+ epsrox = 3.9
+ toxe = 3E-9
+ toxp = 2.8E-9
+ toxm = 3E-9
+ xj = 1E-7
* + gamma1 = 1.2
* + gamma2 = 0.2
+ ndep = 1.7E17
* + nsub = 6E16
+ ngate = 1E23
+ nsd = 1E20
* + vbx = -42
* + xt = 1.55E-7
+ rsh = 0
+ rshg = 0.1
+ phin = 0
+ wint = 0
+ wl = 0
+ wln = 1
+ ww = 0
+ wwn = 1
+ wwl = 0
+ lint = 0
+ ll = 0
+ lln = 1
+ lw = 0
+ lwn = 1
+ lwl = 0
+ llc = 0
+ lwc = 0
+ lwlc = 0
+ wlc = 0
+ wwc = 0
+ wwlc = 0
+ dwg = 0
+ dwb = 0
+ xl = 0
+ xw = 0
+ dmcg = 0
+ dmci = 0
+ dmdg = 0
+ dmcgt = 0
+ dwj = 0
+ xgw = 0
+ xgl = 0
+ ngcon = 1
+ vth0 = 0.5
+ vfb = -1
+ k1 = 0.5
+ k2 = -0.0186
+ k3 = 0
+ k3b = 0
+ w0 = 1E-7
+ lpe0 = 1.74E-7
+ lpeb = 0
+ vbm = -3
+ dvtp0 = 5E-7
+ dvtp1 = 0
+ dvt0 = 2.2
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = 0
+ dvt1w = 5.3
+ dvt2w = -0.032
+ vfbsdoff = 0
+ u0 = 0.05
+ ua = 1E-9
+ ub = 1E-18
+ uc = -4.65E-11
+ ud = 0
+ up = 0
+ lp = 1E-7
+ eu = 1.67
+ vsat = 8E4
+ a0 = 1
+ ags = 0
+ b0 = 0
+ b1 = 0
+ keta = -0.047
+ a1 = 0
+ a2 = 1
+ rdsw = 200
+ rdswmin = 0
+ rdw = 100
+ rdwmin = 0
+ rsw = 100
+ rswmin = 0
+ prwb = 0
+ prwg = 0
+ wr = 1
+ voff = -0.08
+ voffl = 0
+ minv = 0
+ nfactor = 1
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
+ cit = 0
+ cdsc = 2.4E-4
+ cdscb = 0
+ cdscd = 0
+ pclm = 0.5
+ pdiblc1 = 0.39
+ pdiblc2 = 8.6E-3
+ pdiblcb = 0
+ drout = 0.56
+ pscbe1 = 5E9
+ pscbe2 = 5E-6
+ pvag = 0
+ delta = 0.01
+ fprout = 0
+ pdits = 1E-3
+ pditsl = 1
+ pditsd = 0
+ lambda = 0
+ vtl = 0
+ lc = 0
+ xn = 3
+ alpha0 = 0
+ alpha1 = 0
+ beta0 = 15
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1
+ aigbinv = 0.05
+ bigbinv = 0
+ cigbinv = 6E-3
+ eigbinv = 1.1
+ nigbinv = 3
+ aigc = 0.054
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 5E-9
+ nigc = 1
+ poxedge = 1
+ pigcd = 1
+ ntox = 1
+ toxref = 3E-9
+ agidl = 0
+ bgidl = 2.3E9
+ cgidl = 0.5
+ egidl = 0.8
+ xpart = 0
+ cgso = 5E-11
+ cgdo = 5E-11
+ cgbo = 1E-12
+ ckappas = 0.6
+ ckappad = 0.6
+ cf = 5E-11
+ clc = 1E-7
+ cle = 0.6
+ dlc = 0
+ dwc = 0
+ vfbcv = -1
+ noff = 1
+ voffcv = 0
+ acde = 1
+ moin = 15
+ cgsl = 1E-10
+ cgdl = 1E-10
+ ijthsrev = 0.1
+ ijthdrev = 0.1
+ ijthsfwd = 0.1
+ ijthdfwd = 0.1
+ xjbvs = 1
+ xjbvd = 1
+ bvs = 10
+ bvd = 10
+ jss = 1E-4
+ jsd = 1E-4
+ jsws = 1E-14
+ jswd = 1E-14
+ jswgs = 1E-13
+ jswgd = 1E-14
+ jtss = 0
+ jtsd = 0
+ jtssws = 0
+ jtsswd = 0
+ jtsswgs = 0
+ jtsswgd = 0
+ njts = 20
+ njtssw = 20
+ njtsswg = 20
+ xtss = 0.02
+ xtsd = 0.02
+ xtssws = 0.02
+ xtsswd = 0.02
+ xtsswgs = 0.02
+ xtsswgd = 0.02
+ vtss = 10
+ vtsd = 10
+ vtssws = 10
+ vtsswd = 10
+ vtsswgs = 10
+ vtsswgd = 10
+ tnjts = 0
+ tnjtssw = 0
+ tnjtsswg = 0
+ cjs = 5E-4
+ cjd = 5E-4
+ mjs = 0.5
+ mjd = 0.5
+ mjsws = 0.33
+ mjswd = 0.33
+ cjsws = 1E-10
+ cjswd = 1E-10
+ cjswgs = 5E-10
+ cjswgd = 5E-10
+ mjswgs = 0.33
+ mjswgd = 0.33
+ pbs = 0.8
+ pbd = 0.8
+ pbsws = 0.8
+ pbswd = 0.8
+ pbswgs = 0.8
+ pbswgd = 0.8
+ tnom = 25
+ ute = -1.5
+ kt1 = -0.11
+ kt1l = 0
+ kt2 = 0.022
+ ua1 = 6.71E-3
+ ub1 = -3.35E-3
+ uc1 = 4.1E-3
+ ud1 = 0
+ at = 8.13E-3
+ prt = 0
+ njs = 1
+ njd = 1
+ xtis = 3
+ xtid = 3
+ tpb = 0
+ tpbsw = 0
+ tpbswg = 0
+ tcj = 0
+ tcjsw = 0
+ tcjswg = 0
+ tvoff = 0
+ tvfbsdoff = 0
+ saref = 1E-6
+ sbref = 1E-6
+ wlod = 0
+ ku0 = 0
+ kvsat = 0
+ kvth0 = 0
+ tku0 = 0
+ llodku0 = 1
+ wlodku0 = 1
+ llodvth = 1
+ wlodvth = 1
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0
+ lkvth0 = 0
+ wkvth0 = 0
+ pkvth0 = 0
+ stk2 = 0
+ lodk2 = 1
+ steta0 = 0
+ lodeta0 = 1
+ web = 0
+ wec = 0
+ kvth0we = 0
+ k2we = 0
+ ku0we = 0
+ scref = 1E-6
+ wmin = 0.28E-6
+ lmin = 0.22E-6
+ bin_pvsat = 0
+ bin_prdsw = 0
+ bin_ppclm = 0
+ bin_wketa = 0
+ bin_lketa = 0
+ bin_pketa = 0
+ bin_wk3 = 0
+ bin_wk3b = 0

.model nch nmos version=4.8 level=54
* model parameters
+ binunit = 'binunit'
+ paramchk = 'paramchk'
+ mobmod = 'mobmod'
+ capmod = 'capmod'
+ rdsmod = 'rdsmod'
+ igcmod = 'igcmod'
+ igbmod = 'igbmod'
+ rbodymod = 'rbodymod'
+ trnqsmod = 'trnqsmod'
+ acnqsmod = 'acnqsmod'
+ fnoimod = 'fnoimod'
+ tnoimod = 'tnoimod'
+ diomod = 'diomod'
+ tempmod = 'tempmod'
+ permod = 'permod'
+ geomod = 'geomod'
+ rgeomod = 'rgeomod'
+ rgatemod = 'rgatemod'
+ wpemod = 'wpemod'
+ lmin = 'lmin'
+ lmax = 'lmax'
+ wmin = 'wmin'
+ wmax = 'wmax'
+ epsrox = 'epsrox'
+ toxe = 'toxe'
+ toxp = 'toxp'
+ toxm = 'toxm'
+ xj = 'xj'
* + gamma1 = 'gamma1'
* + gamma2 = 'gamma2'
+ ndep = 'ndep'
* + nsub = 'nsub'
+ ngate = 'ngate'
+ nsd = 'nsd'
* + vbx = 'vbx'
* + xt = 'xt'
+ rsh = 'rsh'
+ rshg = 'rshg'
+ phin = 'phin'
+ wint = 'wint'
+ wl = 'wl'
+ wln = 'wln'
+ ww = 'ww'
+ wwn = 'wwn'
+ wwl = 'wwl'
+ lint = 'lint'
+ ll = 'll'
+ lln = 'lln'
+ lw = 'lw'
+ lwn = 'lwn'
+ lwl = 'lwl'
+ llc = 'llc'
+ lwc = 'lwc'
+ lwlc = 'lwlc'
+ wlc = 'wlc'
+ wwc = 'wwc'
+ wwlc = 'wwlc'
+ dwg = 'dwg'
+ dwb = 'dwb'
+ xl = 'xl'
+ xw = 'xw'
+ dmcg = 'dmcg'
+ dmci = 'dmci'
+ dmdg = 'dmdg'
+ dmcgt = 'dmcgt'
+ dwj = 'dwj'
+ xgw = 'xgw'
+ xgl = 'xgl'
+ ngcon = 'ngcon'
+ vth0 = 'vth0'
+ vfb = 'vfb'
+ k1 = 'k1'
+ k2 = 'k2'
+ w0 = 'w0'
+ lpe0 = 'lpe0'
+ lpeb = 'lpeb'
+ vbm = 'vbm'
+ dvtp0 = 'dvtp0'
+ dvtp1 = 'dvtp1'
+ dvt0 = 'dvt0'
+ dvt1 = 'dvt1'
+ dvt2 = 'dvt2'
+ dvt0w = 'dvt0w'
+ dvt1w = 'dvt1w'
+ dvt2w = 'dvt2w'
+ vfbsdoff = 'vfbsdoff'
+ u0 = 'u0'
+ ua = 'ua'
+ ub = 'ub'
+ uc = 'uc'
+ ud = 'ud'
+ up = 'up'
+ lp = 'lp'
+ eu = 'eu'
+ a0 = 'a0'
+ ags = 'ags'
+ b0 = 'b0'
+ b1 = 'b1'
+ a1 = 'a1'
+ a2 = 'a2'
+ rdw = 'rdw'
+ rdswmin = 'rdswmin'
+ rdwmin = 'rdwmin'
+ rsw = 'rsw'
+ rswmin = 'rswmin'
+ prwb = 'prwb'
+ prwg = 'prwg'
+ wr = 'wr'
+ voff = 'voff'
+ voffl = 'voffl'
+ minv = 'minv'
+ nfactor = 'nfactor'
+ eta0 = 'eta0'
+ etab = 'etab'
+ dsub = 'dsub'
+ cit = 'cit'
+ cdsc = 'cdsc'
+ cdscb = 'cdscb'
+ cdscd = 'cdscd'
+ pdiblc1 = 'pdiblc1'
+ pdiblc2 = 'pdiblc2'
+ pdiblcb = 'pdiblcb'
+ drout = 'drout'
+ pscbe1 = 'pscbe1'
+ pscbe2 = 'pscbe2'
+ pvag = 'pvag'
+ delta = 'delta'
+ fprout = 'fprout'
+ pdits = 'pdits'
+ pditsl = 'pditsl'
+ pditsd = 'pditsd'
+ lambda = 'lambda'
+ vtl = 'vtl'
+ lc = 'lc'
+ xn = 'xn'
+ alpha0 = 'alpha0'
+ alpha1 = 'alpha1'
+ beta0 = 'beta0'
+ aigbacc = 'aigbacc'
+ bigbacc = 'bigbacc'
+ cigbacc = 'cigbacc'
+ nigbacc = 'nigbacc'
+ aigbinv = 'aigbinv'
+ bigbinv = 'bigbinv'
+ cigbinv = 'cigbinv'
+ eigbinv = 'eigbinv'
+ nigbinv = 'nigbinv'
+ aigc = 'aigc'
+ bigc = 'bigc'
+ cigc = 'cigc'
+ aigsd = 'aigsd'
+ bigsd = 'bigsd'
+ cigsd = 'cigsd'
+ dlcig = 'dlcig'
+ nigc = 'nigc'
+ poxedge = 'poxedge'
+ pigcd = 'pigcd'
+ ntox = 'ntox'
+ toxref = 'toxref'
+ agidl = 'agidl'
+ bgidl = 'bgidl'
+ cgidl = 'cgidl'
+ egidl = 'egidl'
+ xpart = 'xpart'
+ cgso = 'cgso'
+ cgdo = 'cgdo'
+ cgbo = 'cgbo'
+ ckappas = 'ckappas'
+ ckappad = 'ckappad'
+ cf = 'cf'
+ clc = 'clc'
+ cle = 'cle'
+ dlc = 'dlc'
+ dwc = 'dwc'
+ vfbcv = 'vfbcv'
+ noff = 'noff'
+ voffcv = 'voffcv'
+ acde = 'acde'
+ moin = 'moin'
+ cgsl = 'cgsl'
+ cgdl = 'cgdl'
+ ijthsrev = 'ijthsrev'
+ ijthdrev = 'ijthdrev'
+ ijthsfwd = 'ijthsfwd'
+ ijthdfwd = 'ijthdfwd'
+ xjbvs = 'xjbvs'
+ xjbvd = 'xjbvd'
+ bvs = 'bvs'
+ bvd = 'bvd'
+ jss = 'jss'
+ jsd = 'jsd'
+ jsws = 'jsws'
+ jswd = 'jswd'
+ jswgs = 'jswgs'
+ jswgd = 'jswgd'
+ jtss = 'jtss'
+ jtsd = 'jtsd'
+ jtssws = 'jtssws'
+ jtsswd = 'jtsswd'
+ jtsswgs = 'jtsswgs'
+ jtsswgd = 'jtsswgd'
+ njts = 'njts'
+ njtssw = 'njtssw'
+ njtsswg = 'njtsswg'
+ xtss = 'xtss'
+ xtsd = 'xtsd'
+ xtssws = 'xtssws'
+ xtsswd = 'xtsswd'
+ xtsswgs = 'xtsswgs'
+ xtsswgd = 'xtsswgd'
+ vtss = 'vtss'
+ vtsd = 'vtsd'
+ vtssws = 'vtssws'
+ vtsswd = 'vtsswd'
+ vtsswgs = 'vtsswgs'
+ vtsswgd = 'vtsswgd'
+ tnjts = 'tnjts'
+ tnjtssw = 'tnjtssw'
+ tnjtsswg = 'tnjtsswg'
+ cjs = 'cjs'
+ cjd = 'cjd'
+ mjs = 'mjs'
+ mjd = 'mjd'
+ mjsws = 'mjsws'
+ mjswd = 'mjswd'
+ cjsws = 'cjsws'
+ cjswd = 'cjswd'
+ cjswgs = 'cjswgs'
+ cjswgd = 'cjswgd'
+ mjswgs = 'mjswgs'
+ mjswgd = 'mjswgd'
+ pbs = 'pbs'
+ pbd = 'pbd'
+ pbsws = 'pbsws'
+ pbswd = 'pbswd'
+ pbswgs = 'pbswgs'
+ pbswgd = 'pbswgd'
+ tnom = 'tnom'
+ ute = 'ute'
+ kt1 = 'kt1'
+ kt1l = 'kt1l'
+ kt2 = 'kt2'
+ ua1 = 'ua1'
+ ub1 = 'ub1'
+ uc1 = 'uc1'
+ ud1 = 'ud1'
+ at = 'at'
+ prt = 'prt'
+ njs = 'njs'
+ njd = 'njd'
+ xtis = 'xtis'
+ xtid = 'xtid'
+ tpb = 'tpb'
+ tpbsw = 'tpbsw'
+ tpbswg = 'tpbswg'
+ tcj = 'tcj'
+ tcjsw = 'tcjsw'
+ tcjswg = 'tcjswg'
+ tvoff = 'tvoff'
+ tvfbsdoff = 'tvfbsdoff'
+ saref = 'saref'
+ sbref = 'sbref'
+ wlod = 'wlod'
+ ku0 = 'ku0'
+ kvsat = 'kvsat'
+ kvth0 = 'kvth0'
+ tku0 = 'tku0'
+ llodku0 = 'llodku0'
+ wlodku0 = 'wlodku0'
+ llodvth = 'llodvth'
+ wlodvth = 'wlodvth'
+ lku0 = 'lku0'
+ wku0 = 'wku0'
+ pku0 = 'pku0'
+ lkvth0 = 'lkvth0'
+ wkvth0 = 'wkvth0'
+ pkvth0 = 'pkvth0'
+ stk2 = 'stk2'
+ lodk2 = 'lodk2'
+ steta0 = 'steta0'
+ lodeta0 = 'lodeta0'
+ web = 'web'
+ wec = 'wec'
+ kvth0we = 'kvth0we'
+ k2we = 'k2we'
+ ku0we = 'ku0we'
+ scref = 'scref'
+ vsat = 'vsat'
+ pvsat = 'vsat * bin_pvsat * (lmin * wmin)'
+ rdsw = 'rdsw'
+ prdsw = 'rdsw * bin_prdsw * (lmin * wmin)'
+ pclm = 'pclm'
+ ppclm = 'pclm * bin_ppclm * (lmin * wmin)'
+ keta = 'keta'
+ lketa = 'keta * bin_lketa * lmin'
+ wketa = 'keta * bin_wketa * wmin'
+ pketa = 'keta * bin_pketa * (lmin * wmin)'
+ k3 = 'k3'
+ wk3 = 'k3 * bin_wk3 * wmin'
+ k3b = 'k3b'
+ wk3b = 'k3b * bin_wk3b * wmin'


m1 d g s b nch
+ l = l
+ w = w
+ nf = nf
+ m = m
+ sa = sa
+ sb = sb
+ sc = sc
+ sca = sca
+ scb = scb
+ scc = scc
+ ad = ad
+ pd = pd
+ as = as
+ ps = ps
+ nrs = nrs
+ nrd = nrd

.include dut1.cir

.ends